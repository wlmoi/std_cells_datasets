magic
tech sky130A
timestamp 1745128165
<< locali >>
rect 3715 1440 3800 1455
rect 3715 1435 3730 1440
rect 2230 1410 3730 1435
rect 1320 1365 1345 1400
rect 3715 1385 3730 1410
rect 3790 1385 3800 1440
rect 3715 1370 3800 1385
rect 1300 1350 1360 1365
rect 1300 1320 1315 1350
rect 1345 1320 1360 1350
rect 1300 1305 1360 1320
rect 5640 1210 5715 1225
rect 5640 1185 5650 1210
rect 5700 1185 5715 1210
rect 5640 1165 5715 1185
rect 5650 1120 5670 1165
rect 130 670 150 725
rect 3420 710 3480 720
rect 3420 703 3425 710
rect 3285 673 3425 703
rect 90 655 160 670
rect 90 615 110 655
rect 145 615 160 655
rect 3420 660 3425 673
rect 3470 703 3480 710
rect 3662 703 3702 837
rect 3470 673 3702 703
rect 3470 660 3480 673
rect 3420 650 3480 660
rect 5560 620 5580 655
rect 90 605 160 615
rect 5550 610 5610 620
rect 5550 575 5560 610
rect 5600 575 5610 610
rect 5550 560 5610 575
rect 3885 475 3960 490
rect 3885 435 3900 475
rect 3940 460 3960 475
rect 3940 435 3995 460
rect 3400 405 3470 420
rect 3885 415 3960 435
rect 3400 365 3420 405
rect 3455 365 3470 405
rect 3400 350 3470 365
rect 645 325 705 340
rect 645 290 660 325
rect 695 320 705 325
rect 695 295 735 320
rect 695 290 705 295
rect 645 265 705 290
<< viali >>
rect 3730 1385 3790 1440
rect 1315 1320 1345 1350
rect 5650 1185 5700 1210
rect 110 615 145 655
rect 3425 660 3470 710
rect 5560 575 5600 610
rect 3900 435 3940 475
rect 3420 365 3455 405
rect 660 290 695 325
<< metal1 >>
rect 3715 1440 3800 1455
rect 3715 1385 3730 1440
rect 3790 1395 3990 1440
rect 3790 1385 3800 1395
rect 3715 1370 3800 1385
rect 1300 1350 1360 1365
rect 1300 1320 1315 1350
rect 1345 1320 1360 1350
rect 1300 1305 1360 1320
rect 5640 1210 5715 1225
rect 5640 1185 5650 1210
rect 5700 1185 5715 1210
rect 5640 1165 5715 1185
rect 3420 710 3480 720
rect 90 655 160 670
rect 90 615 110 655
rect 145 615 160 655
rect 3420 660 3425 710
rect 3470 660 3480 710
rect 3420 650 3480 660
rect 3795 650 3930 675
rect 90 605 160 615
rect 2940 435 2950 455
rect 2925 410 2950 435
rect 3400 410 3470 420
rect 3795 410 3820 650
rect 5550 610 5610 620
rect 5550 575 5560 610
rect 5600 575 5610 610
rect 5550 560 5610 575
rect 3885 475 3960 490
rect 3885 435 3900 475
rect 3940 435 3960 475
rect 3885 415 3960 435
rect 2925 405 3820 410
rect 2925 380 3420 405
rect 3400 365 3420 380
rect 3455 380 3820 405
rect 3455 365 3470 380
rect 3400 350 3470 365
rect 645 325 705 340
rect 645 290 660 325
rect 695 290 705 325
rect 645 265 705 290
use ff_common  ff_common_0
timestamp 1744728648
transform 1 0 3841 0 1 640
box -210 -535 1975 825
use mux_common  mux_common_0
timestamp 1744708989
transform 1 0 265 0 1 515
box -265 -515 3020 1219
<< labels >>
rlabel viali 110 615 145 655 1 in_sel
rlabel viali 660 290 695 325 1 in_b
rlabel viali 3420 365 3455 405 1 gnd
rlabel viali 3730 1385 3790 1440 1 vdd
rlabel viali 5650 1185 5700 1210 1 out_q
rlabel viali 5560 575 5600 610 1 out_q_not
rlabel viali 3900 435 3940 475 1 in_clk
rlabel viali 3425 660 3470 710 1 out_mux
rlabel viali 1315 1320 1345 1350 1 in_a
<< end >>
