magic
tech sky130A
timestamp 1744191774
<< nwell >>
rect -225 -20 55 105
rect 240 -20 515 105
<< nmos >>
rect -45 -165 -30 -100
rect 330 -165 345 -100
<< pmos >>
rect -45 5 -30 70
rect 330 5 345 70
<< ndiff >>
rect -100 -115 -45 -100
rect -100 -150 -85 -115
rect -65 -150 -45 -115
rect -100 -165 -45 -150
rect -30 -115 20 -100
rect -30 -150 -10 -115
rect 10 -150 20 -115
rect -30 -165 20 -150
rect 280 -115 330 -100
rect 280 -155 290 -115
rect 310 -155 330 -115
rect 280 -165 330 -155
rect 345 -115 400 -100
rect 345 -155 365 -115
rect 385 -155 400 -115
rect 345 -165 400 -155
<< pdiff >>
rect -95 55 -45 70
rect -95 20 -85 55
rect -65 20 -45 55
rect -95 5 -45 20
rect -30 55 20 70
rect -30 20 -10 55
rect 10 20 20 55
rect -30 5 20 20
rect 275 55 330 70
rect 275 15 285 55
rect 310 15 330 55
rect 275 5 330 15
rect 345 55 400 70
rect 345 15 365 55
rect 390 15 400 55
rect 345 5 400 15
<< ndiffc >>
rect -85 -150 -65 -115
rect -10 -150 10 -115
rect 290 -155 310 -115
rect 365 -155 385 -115
<< pdiffc >>
rect -85 20 -65 55
rect -10 20 10 55
rect 285 15 310 55
rect 365 15 390 55
<< psubdiff >>
rect 245 -230 320 -210
rect 245 -260 265 -230
rect 300 -260 320 -230
rect 245 -275 320 -260
<< nsubdiff >>
rect -190 50 -130 70
rect -190 25 -170 50
rect -150 25 -130 50
rect -190 5 -130 25
rect 440 55 485 70
rect 440 20 450 55
rect 475 20 485 55
rect 440 5 485 20
<< psubdiffcont >>
rect 265 -260 300 -230
<< nsubdiffcont >>
rect -170 25 -150 50
rect 450 20 475 55
<< poly >>
rect -45 70 -30 85
rect 330 70 345 85
rect -45 -40 -30 5
rect -85 -50 -30 -40
rect -85 -75 -75 -50
rect -55 -75 -30 -50
rect -85 -80 -30 -75
rect -45 -100 -30 -80
rect 330 -35 345 5
rect 330 -45 390 -35
rect 330 -70 355 -45
rect 380 -70 390 -45
rect 330 -80 390 -70
rect 330 -100 345 -80
rect -45 -180 -30 -165
rect 330 -180 345 -165
<< polycont >>
rect -75 -75 -55 -50
rect 355 -70 380 -45
<< locali >>
rect 135 175 620 200
rect -190 50 -130 70
rect -95 55 -55 70
rect -95 50 -85 55
rect -190 25 -170 50
rect -150 25 -85 50
rect -190 5 -130 25
rect -95 20 -85 25
rect -65 20 -55 55
rect -95 5 -55 20
rect -20 55 20 70
rect -20 20 -10 55
rect 10 20 20 55
rect -20 5 20 20
rect -85 -50 -45 -40
rect -85 -75 -75 -50
rect -55 -75 -45 -50
rect -85 -80 -45 -75
rect -10 -50 10 5
rect 135 -50 160 175
rect 275 55 320 70
rect 275 15 285 55
rect 310 15 320 55
rect 275 5 320 15
rect 355 55 400 70
rect 355 15 365 55
rect 390 50 400 55
rect 440 55 485 70
rect 440 50 450 55
rect 390 30 450 50
rect 390 15 400 30
rect 355 5 400 15
rect 440 20 450 30
rect 475 20 485 55
rect 440 5 485 20
rect 290 -50 310 5
rect -10 -70 310 -50
rect 345 -45 390 -35
rect 345 -70 355 -45
rect 380 -70 390 -45
rect -10 -100 10 -70
rect 345 -80 390 -70
rect 595 -100 620 175
rect -100 -115 -55 -100
rect -100 -150 -85 -115
rect -65 -150 -55 -115
rect -100 -165 -55 -150
rect -20 -115 20 -100
rect -20 -150 -10 -115
rect 10 -150 20 -115
rect -20 -165 20 -150
rect 280 -115 320 -100
rect 280 -155 290 -115
rect 310 -155 320 -115
rect 280 -165 320 -155
rect 355 -115 400 -100
rect 355 -155 365 -115
rect 385 -155 400 -115
rect 595 -125 675 -100
rect 355 -165 400 -155
rect -85 -325 -65 -165
rect 290 -210 310 -165
rect 245 -230 320 -210
rect 245 -260 265 -230
rect 300 -260 320 -230
rect 245 -275 320 -260
rect 370 -325 390 -165
rect -85 -345 390 -325
<< viali >>
rect -170 25 -150 50
rect 450 20 475 55
rect 265 -260 300 -230
<< metal1 >>
rect -190 50 -130 70
rect -190 25 -170 50
rect -150 25 -130 50
rect -190 5 -130 25
rect 440 55 485 70
rect 440 20 450 55
rect 475 20 485 55
rect 440 5 485 20
rect 245 -230 320 -210
rect 245 -260 265 -230
rect 300 -260 320 -230
rect 245 -275 320 -260
use inv2  inv2_0 /foss/designs/eda/inverter
timestamp 1743223184
transform 1 0 815 0 1 -10
box -140 -335 125 175
<< labels >>
rlabel polycont -75 -75 -55 -50 1 in1
rlabel nwell -170 25 -150 50 1 vcc
rlabel polycont 355 -70 380 -45 1 in2
rlabel metal1 265 -260 300 -230 1 gnd
rlabel nwell 450 20 475 55 1 vcc
rlabel space 845 -125 870 -100 1 out
rlabel space 800 100 840 130 1 vcc
rlabel space 815 -330 840 -310 1 gnd
<< end >>
