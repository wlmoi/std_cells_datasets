magic
tech sky130A
timestamp 1744185391
<< nwell >>
rect -225 -20 315 105
<< nmos >>
rect -45 -165 -30 -100
rect 130 -165 145 -100
<< pmos >>
rect -45 5 -30 70
rect 130 5 145 70
<< ndiff >>
rect -100 -115 -45 -100
rect -100 -150 -85 -115
rect -65 -150 -45 -115
rect -100 -165 -45 -150
rect -30 -115 20 -100
rect -30 -150 -10 -115
rect 10 -150 20 -115
rect -30 -165 20 -150
rect 80 -115 130 -100
rect 80 -155 90 -115
rect 110 -155 130 -115
rect 80 -165 130 -155
rect 145 -115 200 -100
rect 145 -155 165 -115
rect 185 -155 200 -115
rect 145 -165 200 -155
<< pdiff >>
rect -95 55 -45 70
rect -95 20 -85 55
rect -65 20 -45 55
rect -95 5 -45 20
rect -30 55 20 70
rect -30 20 -10 55
rect 10 20 20 55
rect -30 5 20 20
rect 75 55 130 70
rect 75 15 85 55
rect 110 15 130 55
rect 75 5 130 15
rect 145 55 200 70
rect 145 15 165 55
rect 190 15 200 55
rect 145 5 200 15
<< ndiffc >>
rect -85 -150 -65 -115
rect -10 -150 10 -115
rect 90 -155 110 -115
rect 165 -155 185 -115
<< pdiffc >>
rect -85 20 -65 55
rect -10 20 10 55
rect 85 15 110 55
rect 165 15 190 55
<< psubdiff >>
rect 45 -230 120 -210
rect 45 -260 65 -230
rect 100 -260 120 -230
rect 45 -275 120 -260
<< nsubdiff >>
rect -190 50 -130 70
rect -190 25 -170 50
rect -150 25 -130 50
rect -190 5 -130 25
rect 240 55 285 70
rect 240 20 250 55
rect 275 20 285 55
rect 240 5 285 20
<< psubdiffcont >>
rect 65 -260 100 -230
<< nsubdiffcont >>
rect -170 25 -150 50
rect 250 20 275 55
<< poly >>
rect -45 70 -30 85
rect 130 70 145 85
rect -45 -40 -30 5
rect -85 -50 -30 -40
rect -85 -75 -75 -50
rect -55 -75 -30 -50
rect -85 -80 -30 -75
rect -45 -100 -30 -80
rect 130 -35 145 5
rect 130 -45 190 -35
rect 130 -70 155 -45
rect 180 -70 190 -45
rect 130 -80 190 -70
rect 130 -100 145 -80
rect -45 -180 -30 -165
rect 130 -180 145 -165
<< polycont >>
rect -75 -75 -55 -50
rect 155 -70 180 -45
<< locali >>
rect -190 50 -130 70
rect -95 55 -55 70
rect -95 50 -85 55
rect -190 25 -170 50
rect -150 25 -85 50
rect -190 5 -130 25
rect -95 20 -85 25
rect -65 20 -55 55
rect -95 5 -55 20
rect -20 55 20 70
rect -20 20 -10 55
rect 10 20 20 55
rect -20 5 20 20
rect 75 55 120 70
rect 75 15 85 55
rect 110 15 120 55
rect 75 5 120 15
rect 155 55 200 70
rect 155 15 165 55
rect 190 50 200 55
rect 240 55 285 70
rect 240 50 250 55
rect 190 30 250 50
rect 190 15 200 30
rect 155 5 200 15
rect 240 20 250 30
rect 275 20 285 55
rect 240 5 285 20
rect -10 -35 10 5
rect 90 -35 110 5
rect -10 -40 110 -35
rect -85 -50 -45 -40
rect -85 -75 -75 -50
rect -55 -75 -45 -50
rect -85 -80 -45 -75
rect -10 -65 25 -40
rect 60 -65 110 -40
rect -10 -70 110 -65
rect 145 -45 190 -35
rect 145 -70 155 -45
rect 180 -70 190 -45
rect -10 -100 10 -70
rect 145 -80 190 -70
rect -100 -115 -55 -100
rect -100 -150 -85 -115
rect -65 -150 -55 -115
rect -100 -165 -55 -150
rect -20 -115 20 -100
rect -20 -150 -10 -115
rect 10 -150 20 -115
rect -20 -165 20 -150
rect 80 -115 120 -100
rect 80 -155 90 -115
rect 110 -155 120 -115
rect 80 -165 120 -155
rect 155 -115 200 -100
rect 155 -155 165 -115
rect 185 -155 200 -115
rect 155 -165 200 -155
rect -85 -325 -65 -165
rect 90 -210 110 -165
rect 45 -230 120 -210
rect 45 -260 65 -230
rect 100 -260 120 -230
rect 45 -275 120 -260
rect 170 -325 190 -165
rect -85 -345 190 -325
<< viali >>
rect -170 25 -150 50
rect 250 20 275 55
rect 25 -65 60 -40
rect 65 -260 100 -230
<< metal1 >>
rect -190 50 -130 70
rect -190 25 -170 50
rect -150 25 -130 50
rect -190 5 -130 25
rect 240 55 285 70
rect 240 20 250 55
rect 275 20 285 55
rect 240 5 285 20
rect -10 -40 110 -35
rect -10 -65 25 -40
rect 60 -65 110 -40
rect -10 -70 110 -65
rect 45 -230 120 -210
rect 45 -260 65 -230
rect 100 -260 120 -230
rect 45 -275 120 -260
<< labels >>
rlabel polycont -75 -75 -55 -50 1 in1
rlabel polycont 155 -70 180 -45 1 in2
rlabel metal1 65 -260 100 -230 1 gnd
rlabel nwell -170 25 -150 50 1 vcc
rlabel nwell 250 20 275 55 1 vcc
rlabel viali 25 -65 60 -40 1 out
<< end >>
