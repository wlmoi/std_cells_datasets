magic
tech sky130A
timestamp 1744814206
<< locali >>
rect 1035 810 1120 825
rect 1035 770 1055 810
rect 1105 770 1120 810
rect 1035 760 1120 770
rect 495 580 555 590
rect 915 585 970 595
rect 1215 585 1260 595
rect 1630 585 1690 595
rect 495 575 505 580
rect -70 555 505 575
rect 540 560 595 580
rect 870 560 925 585
rect 540 555 555 560
rect -210 255 -115 270
rect -210 205 -200 255
rect -130 250 -115 255
rect -70 250 -45 555
rect 495 540 555 555
rect 915 550 925 560
rect 960 565 1015 585
rect 960 550 970 565
rect 915 540 970 550
rect 900 460 950 470
rect 900 440 910 460
rect 940 440 950 460
rect 900 425 950 440
rect -130 220 0 250
rect 275 245 335 255
rect 205 225 285 245
rect 275 220 285 225
rect 320 220 335 245
rect -130 205 -115 220
rect 275 210 335 220
rect -210 190 -115 205
rect 150 -170 230 -150
rect 150 -210 165 -170
rect 215 -210 230 -170
rect 150 -230 230 -210
rect 185 -460 215 -230
rect 300 -410 325 210
rect 995 60 1015 565
rect 1215 555 1225 585
rect 1250 560 1300 585
rect 1575 580 1690 585
rect 1250 555 1260 560
rect 1575 555 1640 580
rect 1680 560 1735 580
rect 1680 555 1690 560
rect 1215 550 1260 555
rect 1630 545 1690 555
rect 1045 260 1125 280
rect 1045 225 1065 260
rect 1105 225 1125 260
rect 1045 205 1125 225
rect 1165 235 1655 260
rect 1165 155 1190 235
rect 1140 145 1210 155
rect 1140 110 1150 145
rect 1200 110 1210 145
rect 1140 100 1210 110
rect 905 45 955 55
rect 905 15 915 45
rect 945 15 955 45
rect 995 40 1140 60
rect 905 10 955 15
rect 495 -60 545 -50
rect 495 -85 505 -60
rect 535 -85 545 -60
rect 910 -70 970 -60
rect 910 -75 920 -70
rect 495 -95 545 -85
rect 865 -100 920 -75
rect 960 -75 970 -70
rect 960 -100 1085 -75
rect 910 -110 970 -100
rect 995 -205 1040 -195
rect 995 -230 1005 -205
rect 1030 -230 1040 -205
rect 995 -240 1040 -230
rect 1010 -340 1030 -240
rect 960 -355 1030 -340
rect 960 -380 980 -355
rect 1015 -380 1030 -355
rect 960 -390 1030 -380
rect 1060 -410 1085 -100
rect 300 -435 1085 -410
rect 1115 -460 1140 40
rect 1200 -60 1255 -50
rect 1630 -55 1655 235
rect 1710 75 1735 560
rect 1790 475 1885 485
rect 1790 435 1805 475
rect 1875 435 1885 475
rect 1790 420 1885 435
rect 1685 60 1750 75
rect 1685 30 1695 60
rect 1740 30 1750 60
rect 1685 10 1750 30
rect 1200 -90 1215 -60
rect 1245 -70 1255 -60
rect 1615 -65 1665 -55
rect 1615 -70 1625 -65
rect 1245 -90 1300 -70
rect 1575 -90 1625 -70
rect 1655 -90 1665 -65
rect 1200 -100 1255 -90
rect 1615 -100 1665 -90
rect 185 -485 1140 -460
rect 1810 -485 1835 420
rect 1790 -500 1860 -485
rect 1790 -520 1810 -500
rect 1845 -520 1860 -500
rect 1790 -535 1860 -520
<< viali >>
rect 1055 770 1105 810
rect 505 555 540 580
rect -200 205 -130 255
rect 925 550 960 585
rect 910 440 940 460
rect 285 220 320 245
rect 165 -210 215 -170
rect 1225 555 1250 585
rect 1640 555 1680 580
rect 1065 225 1105 260
rect 1150 110 1200 145
rect 915 15 945 45
rect 505 -85 535 -60
rect 920 -100 960 -70
rect 1005 -230 1030 -205
rect 980 -380 1015 -355
rect 1805 435 1875 475
rect 1695 30 1740 60
rect 1215 -90 1245 -60
rect 1625 -90 1655 -65
rect 1810 -520 1845 -500
<< metal1 >>
rect 1035 810 1120 825
rect 1035 800 1055 810
rect 135 775 1055 800
rect 135 770 955 775
rect 135 490 160 770
rect 505 700 530 770
rect 935 700 955 770
rect 1035 770 1055 775
rect 1105 800 1120 810
rect 1105 775 1975 800
rect 1105 770 1120 775
rect 1035 760 1120 770
rect 1215 700 1235 775
rect 1635 700 1655 775
rect 495 580 555 590
rect 495 555 505 580
rect 540 555 555 580
rect 915 585 970 595
rect 495 540 555 555
rect 720 450 740 560
rect 915 550 925 585
rect 960 550 970 585
rect 1215 585 1260 595
rect 1215 555 1225 585
rect 1250 555 1260 585
rect 1630 580 1690 595
rect 1215 550 1260 555
rect 915 540 970 550
rect 900 460 950 470
rect 900 450 910 460
rect 720 440 910 450
rect 940 455 950 460
rect 1230 455 1245 550
rect 940 440 1245 455
rect 1420 460 1445 560
rect 1630 555 1640 580
rect 1680 555 1690 580
rect 1630 545 1690 555
rect 1790 475 1885 485
rect 1790 460 1805 475
rect 1420 440 1805 460
rect 720 435 950 440
rect 900 425 950 435
rect 1790 435 1805 440
rect 1875 435 1885 475
rect 1790 420 1885 435
rect -210 255 -115 270
rect 745 260 775 355
rect 1045 260 1125 280
rect 1460 260 1490 355
rect -210 205 -200 255
rect -130 205 -115 255
rect 275 245 335 255
rect 275 220 285 245
rect 320 220 335 245
rect 275 210 335 220
rect 475 235 1065 260
rect -210 190 -115 205
rect 475 35 500 235
rect 745 130 775 235
rect 1045 225 1065 235
rect 1105 235 1490 260
rect 1105 225 1125 235
rect 1045 205 1125 225
rect 1140 145 1210 155
rect 1140 135 1150 145
rect 920 115 1150 135
rect 920 55 940 115
rect 1140 110 1150 115
rect 1200 110 1210 145
rect 1460 130 1490 235
rect 1140 100 1210 110
rect 1685 60 1750 75
rect 1685 55 1695 60
rect 905 45 955 55
rect 180 10 500 35
rect 715 30 915 45
rect 495 -60 545 -50
rect 495 -65 505 -60
rect 185 -85 505 -65
rect 535 -70 545 -60
rect 535 -85 590 -70
rect 715 -75 730 30
rect 905 15 915 30
rect 945 15 955 45
rect 905 10 955 15
rect 1420 40 1695 55
rect 1200 -60 1255 -50
rect 910 -70 970 -60
rect 185 -150 210 -85
rect 495 -95 590 -85
rect 910 -100 920 -70
rect 960 -100 970 -70
rect 910 -110 970 -100
rect 1020 -85 1215 -60
rect 150 -170 230 -150
rect 150 -210 165 -170
rect 215 -210 230 -170
rect 1020 -195 1040 -85
rect 1200 -90 1215 -85
rect 1245 -90 1255 -60
rect 1420 -70 1440 40
rect 1685 30 1695 40
rect 1740 30 1750 60
rect 1685 10 1750 30
rect 1615 -65 1665 -55
rect 1200 -100 1255 -90
rect 1615 -90 1625 -65
rect 1655 -90 1665 -65
rect 1615 -100 1665 -90
rect 995 -205 1040 -195
rect 150 -230 230 -210
rect 500 -280 530 -215
rect 920 -280 950 -210
rect 995 -230 1005 -205
rect 1030 -230 1040 -205
rect 995 -240 1040 -230
rect 1215 -280 1245 -200
rect 1640 -280 1665 -205
rect 1950 -280 1975 775
rect 500 -315 1975 -280
rect 960 -355 1030 -340
rect 960 -380 980 -355
rect 1015 -380 1030 -355
rect 960 -390 1030 -380
rect 985 -505 1010 -390
rect 1790 -500 1860 -485
rect 1790 -505 1810 -500
rect 985 -520 1810 -505
rect 1845 -520 1860 -500
rect 985 -525 1860 -520
rect 1790 -535 1860 -525
use inverter_common  inverter_common_0
timestamp 1743223184
transform 1 0 140 0 1 335
box -140 -335 125 175
use nand  nand_0
timestamp 1744185391
transform 1 0 680 0 1 630
box -225 -345 315 105
use nand  nand_1
timestamp 1744185391
transform 1 0 675 0 -1 -145
box -225 -345 315 105
use nand  nand_2
timestamp 1744185391
transform 1 0 1385 0 1 630
box -225 -345 315 105
use nand  nand_3
timestamp 1744185391
transform 1 0 1385 0 -1 -140
box -225 -345 315 105
<< labels >>
rlabel viali -200 206 -130 255 1 in_d
rlabel metal1 1065 224 1106 260 1 gnd
rlabel viali 1056 771 1104 810 1 vdd
rlabel metal1 164 -208 214 -169 1 in_clk
rlabel metal1 1805 436 1876 474 1 out_q
rlabel metal1 1695 30 1741 61 1 out_q_not
<< end >>
