magic
tech sky130A
timestamp 1744544585
<< nwell >>
rect -230 -460 -110 85
<< nmos >>
rect -5 -110 65 -90
rect -5 -360 65 -340
<< pmos >>
rect -205 -110 -140 -90
rect -205 -360 -140 -340
<< ndiff >>
rect -5 -40 65 -30
rect -5 -70 10 -40
rect 55 -70 65 -40
rect -5 -90 65 -70
rect -5 -130 65 -110
rect -5 -155 10 -130
rect 50 -155 65 -130
rect -5 -165 65 -155
rect -5 -295 65 -285
rect -5 -320 10 -295
rect 50 -320 65 -295
rect -5 -340 65 -320
rect -5 -380 65 -360
rect -5 -405 10 -380
rect 50 -405 65 -380
rect -5 -415 65 -405
<< pdiff >>
rect -205 -40 -140 -30
rect -205 -70 -195 -40
rect -150 -70 -140 -40
rect -205 -90 -140 -70
rect -205 -130 -140 -110
rect -205 -155 -190 -130
rect -155 -155 -140 -130
rect -205 -165 -140 -155
rect -205 -295 -140 -285
rect -205 -320 -195 -295
rect -150 -320 -140 -295
rect -205 -340 -140 -320
rect -205 -380 -140 -360
rect -205 -405 -195 -380
rect -150 -405 -140 -380
rect -205 -415 -140 -405
<< ndiffc >>
rect 10 -70 55 -40
rect 10 -155 50 -130
rect 10 -320 50 -295
rect 10 -405 50 -380
<< pdiffc >>
rect -195 -70 -150 -40
rect -190 -155 -155 -130
rect -195 -320 -150 -295
rect -195 -405 -150 -380
<< psubdiff >>
rect -5 45 65 60
rect -5 20 15 45
rect 50 20 65 45
rect -5 5 65 20
rect -5 -465 65 -455
rect -5 -495 10 -465
rect 50 -495 65 -465
rect -5 -505 65 -495
<< nsubdiff >>
rect -205 45 -140 60
rect -205 20 -190 45
rect -155 20 -140 45
rect -205 5 -140 20
<< psubdiffcont >>
rect 15 20 50 45
rect 10 -495 50 -465
<< nsubdiffcont >>
rect -190 20 -155 45
<< poly >>
rect -85 -55 -40 -50
rect -85 -85 -75 -55
rect -50 -85 -40 -55
rect -85 -90 -40 -85
rect -220 -110 -205 -90
rect -140 -110 -5 -90
rect 65 -110 80 -90
rect -220 -360 -205 -340
rect -140 -360 -5 -340
rect 65 -360 80 -340
rect -85 -370 -40 -360
rect -85 -395 -75 -370
rect -50 -395 -40 -370
rect -85 -405 -40 -395
<< polycont >>
rect -75 -85 -50 -55
rect -75 -395 -50 -370
<< locali >>
rect -180 105 305 125
rect -180 60 -160 105
rect -205 45 -140 60
rect -205 20 -190 45
rect -155 20 -140 45
rect -205 5 -140 20
rect -5 45 65 60
rect -5 20 15 45
rect 50 25 125 45
rect 50 20 65 25
rect -5 5 65 20
rect -185 -30 -165 5
rect 20 -30 45 5
rect -205 -40 -140 -30
rect -205 -70 -195 -40
rect -150 -70 -140 -40
rect -5 -40 65 -30
rect -205 -80 -140 -70
rect -85 -55 -40 -50
rect -85 -85 -75 -55
rect -50 -85 -40 -55
rect -5 -70 10 -40
rect 55 -70 65 -40
rect -5 -80 65 -70
rect -85 -90 -40 -85
rect -205 -130 -140 -120
rect -5 -130 65 -120
rect -285 -155 -190 -130
rect -155 -155 -140 -130
rect -285 -385 -265 -155
rect -205 -165 -140 -155
rect -85 -155 10 -130
rect 50 -155 65 -130
rect -85 -195 -40 -155
rect -5 -165 65 -155
rect -85 -245 -80 -195
rect -45 -245 -40 -195
rect -205 -295 -140 -285
rect -85 -295 -40 -245
rect -5 -295 65 -285
rect -205 -320 -195 -295
rect -150 -320 10 -295
rect 50 -320 65 -295
rect -205 -330 -140 -320
rect -5 -330 65 -320
rect -85 -370 -40 -360
rect -205 -380 -140 -370
rect -205 -385 -195 -380
rect -285 -405 -195 -385
rect -150 -405 -140 -380
rect -85 -395 -75 -370
rect -50 -395 -40 -370
rect -85 -405 -40 -395
rect -5 -380 65 -370
rect -5 -405 10 -380
rect 50 -405 65 -380
rect -205 -415 -140 -405
rect -5 -415 65 -405
rect 20 -455 40 -415
rect 105 -425 125 25
rect 285 15 305 105
rect 105 -445 230 -425
rect -5 -465 65 -455
rect -5 -495 10 -465
rect 50 -470 65 -465
rect 105 -470 125 -445
rect 50 -490 125 -470
rect 50 -495 65 -490
rect -5 -505 65 -495
<< viali >>
rect -190 20 -155 45
rect 15 20 50 45
rect -80 -245 -45 -195
rect 165 -240 190 -215
rect 10 -495 50 -465
<< metal1 >>
rect -205 45 -140 60
rect -205 20 -190 45
rect -155 20 -140 45
rect -205 5 -140 20
rect -5 45 65 60
rect -5 20 15 45
rect 50 20 65 45
rect -5 5 65 20
rect -85 -195 -40 -130
rect -85 -245 -80 -195
rect -45 -210 -40 -195
rect 150 -210 205 -200
rect -45 -215 205 -210
rect -45 -230 165 -215
rect -45 -245 -40 -230
rect -85 -320 -40 -245
rect 150 -240 165 -230
rect 190 -240 205 -215
rect 150 -255 205 -240
rect -5 -465 65 -455
rect -5 -495 10 -465
rect 50 -495 65 -465
rect -5 -505 65 -495
use inv2  inv2_0 /foss/designs/eda/inverter
timestamp 1743223184
transform 1 0 290 0 1 -125
box -140 -335 125 175
<< labels >>
rlabel metal1 10 -495 50 -465 7 gnd
rlabel metal1 15 20 50 45 7 gnd
rlabel polycont -75 -395 -50 -370 7 in2
rlabel viali -80 -245 -45 -195 7 out
rlabel polycont -75 -85 -50 -55 7 in1
rlabel nwell -190 20 -155 45 7 vdd
<< end >>
