magic
tech sky130A
timestamp 1744220241
<< nwell >>
rect 240 75 430 315
rect -270 -65 430 75
<< nmos >>
rect -30 -235 -10 -155
rect 165 -235 185 -155
rect 350 -360 445 -340
<< pmos >>
rect 285 215 385 235
rect -30 -35 -10 45
rect 165 -35 185 45
<< ndiff >>
rect -100 -170 -30 -155
rect -100 -215 -85 -170
rect -50 -215 -30 -170
rect -100 -235 -30 -215
rect -10 -170 50 -155
rect -10 -215 10 -170
rect 40 -215 50 -170
rect -10 -235 50 -215
rect 100 -170 165 -155
rect 100 -215 115 -170
rect 145 -215 165 -170
rect 100 -235 165 -215
rect 185 -170 245 -155
rect 185 -215 205 -170
rect 235 -215 245 -170
rect 185 -235 245 -215
rect 350 -290 445 -275
rect 350 -320 365 -290
rect 430 -320 445 -290
rect 350 -340 445 -320
rect 350 -385 445 -360
rect 350 -410 365 -385
rect 430 -410 445 -385
rect 350 -425 445 -410
<< pdiff >>
rect 285 280 385 290
rect 285 255 305 280
rect 365 255 385 280
rect 285 235 385 255
rect 285 190 385 215
rect 285 165 305 190
rect 365 165 385 190
rect 285 155 385 165
rect -100 25 -30 45
rect -100 -15 -85 25
rect -55 -15 -30 25
rect -100 -35 -30 -15
rect -10 25 50 45
rect -10 -15 10 25
rect 40 -15 50 25
rect -10 -35 50 -15
rect 100 25 165 45
rect 100 -15 115 25
rect 145 -15 165 25
rect 100 -35 165 -15
rect 185 25 245 45
rect 185 -15 205 25
rect 235 -15 245 25
rect 185 -35 245 -15
<< ndiffc >>
rect -85 -215 -50 -170
rect 10 -215 40 -170
rect 115 -215 145 -170
rect 205 -215 235 -170
rect 365 -320 430 -290
rect 365 -410 430 -385
<< pdiffc >>
rect 305 255 365 280
rect 305 165 365 190
rect -85 -15 -55 25
rect 10 -15 40 25
rect 115 -15 145 25
rect 205 -15 235 25
<< psubdiff >>
rect -220 -175 -145 -155
rect -220 -215 -200 -175
rect -165 -215 -145 -175
rect -220 -235 -145 -215
<< nsubdiff >>
rect -220 25 -145 45
rect -220 -15 -200 25
rect -165 -15 -145 25
rect -220 -35 -145 -15
<< psubdiffcont >>
rect -200 -215 -165 -175
<< nsubdiffcont >>
rect -200 -15 -165 25
<< poly >>
rect 180 245 230 255
rect 180 210 190 245
rect 220 235 230 245
rect 220 215 285 235
rect 385 215 405 235
rect 220 210 230 215
rect 180 200 230 210
rect 165 115 210 125
rect 165 95 175 115
rect 200 95 210 115
rect 165 85 210 95
rect -30 45 -10 60
rect 165 45 185 85
rect -30 -85 -10 -35
rect -80 -95 -10 -85
rect -80 -125 -70 -95
rect -40 -125 -10 -95
rect -80 -135 -10 -125
rect -30 -155 -10 -135
rect 165 -85 185 -35
rect 165 -95 235 -85
rect 165 -125 195 -95
rect 225 -125 235 -95
rect 165 -135 235 -125
rect 165 -155 185 -135
rect -30 -250 -10 -235
rect 165 -265 185 -235
rect 150 -275 200 -265
rect 150 -295 160 -275
rect 190 -295 200 -275
rect 150 -305 200 -295
rect 280 -340 320 -330
rect 280 -360 285 -340
rect 315 -360 350 -340
rect 445 -360 460 -340
rect 280 -370 320 -360
<< polycont >>
rect 190 210 220 245
rect 175 95 200 115
rect -70 -125 -40 -95
rect 195 -125 225 -95
rect 160 -295 190 -275
rect 285 -360 315 -340
<< locali >>
rect 285 280 385 290
rect 285 255 305 280
rect 365 260 580 280
rect 365 255 385 260
rect 180 245 230 255
rect 285 245 385 255
rect 180 235 190 245
rect -330 215 190 235
rect -330 -95 -310 215
rect 115 45 135 215
rect 180 210 190 215
rect 220 210 230 245
rect 180 200 230 210
rect 285 190 385 205
rect 285 175 305 190
rect 180 165 305 175
rect 365 165 385 190
rect 180 155 385 165
rect 180 125 200 155
rect 165 115 210 125
rect 165 95 175 115
rect 200 95 210 115
rect 165 85 210 95
rect -220 25 -145 45
rect -220 -15 -200 25
rect -165 20 -145 25
rect -100 25 -40 45
rect -100 20 -85 25
rect -165 -10 -85 20
rect -165 -15 -145 -10
rect -220 -35 -145 -15
rect -100 -15 -85 -10
rect -55 -15 -40 25
rect -100 -35 -40 -15
rect 0 25 50 45
rect 0 -15 10 25
rect 40 -15 50 25
rect 0 -35 50 -15
rect 100 25 155 45
rect 100 -15 115 25
rect 145 -15 155 25
rect 100 -35 155 -15
rect 195 25 245 45
rect 195 -15 205 25
rect 235 15 245 25
rect 235 -5 320 15
rect 235 -15 245 -5
rect 195 -35 245 -15
rect -80 -95 -30 -85
rect -330 -120 -70 -95
rect -80 -125 -70 -120
rect -40 -125 -30 -95
rect -80 -135 -30 -125
rect 15 -95 35 -35
rect 185 -95 235 -85
rect 15 -115 140 -95
rect 15 -155 35 -115
rect 120 -155 140 -115
rect 185 -125 195 -95
rect 225 -125 235 -95
rect 185 -135 235 -125
rect 300 -120 320 -5
rect 560 -80 580 260
rect 560 -90 630 -80
rect 560 -120 590 -90
rect 300 -125 590 -120
rect 615 -125 630 -90
rect 300 -140 630 -125
rect -220 -175 -145 -155
rect -220 -215 -200 -175
rect -165 -185 -145 -175
rect -100 -170 -40 -155
rect -100 -185 -85 -170
rect -165 -205 -85 -185
rect -165 -215 -145 -205
rect -220 -235 -145 -215
rect -100 -215 -85 -205
rect -50 -215 -40 -170
rect -100 -235 -40 -215
rect 0 -170 50 -155
rect 0 -215 10 -170
rect 40 -215 50 -170
rect 0 -235 50 -215
rect 100 -170 155 -155
rect 100 -215 115 -170
rect 145 -215 155 -170
rect 100 -235 155 -215
rect 195 -170 245 -155
rect 195 -215 205 -170
rect 235 -185 245 -170
rect 300 -185 320 -140
rect 235 -205 320 -185
rect 235 -215 245 -205
rect 195 -235 245 -215
rect 110 -340 130 -235
rect 150 -275 200 -265
rect 150 -295 160 -275
rect 190 -280 200 -275
rect 350 -280 445 -275
rect 190 -290 445 -280
rect 190 -295 365 -290
rect 150 -300 365 -295
rect 150 -305 200 -300
rect 350 -320 365 -300
rect 430 -320 445 -290
rect 350 -330 445 -320
rect 280 -340 320 -330
rect 110 -360 285 -340
rect 315 -360 320 -340
rect 280 -370 320 -360
rect 350 -385 445 -370
rect 560 -385 580 -140
rect 350 -410 365 -385
rect 430 -410 580 -385
rect 350 -425 445 -410
<< viali >>
rect -200 -15 -165 25
rect 590 -125 615 -90
rect -200 -215 -165 -175
<< metal1 >>
rect -220 25 -145 45
rect -220 -15 -200 25
rect -165 -15 -145 25
rect -220 -35 -145 -15
rect 580 -90 630 -80
rect 580 -125 590 -90
rect 615 -125 630 -90
rect 580 -140 630 -125
rect -220 -175 -145 -155
rect -220 -215 -200 -175
rect -165 -215 -145 -175
rect -220 -235 -145 -215
<< labels >>
rlabel nwell -200 -15 -165 25 1 vdd
rlabel metal1 -200 -215 -165 -175 1 gnd
rlabel polycont -70 -125 -40 -95 1 in1
rlabel polycont 195 -125 225 -95 1 in2
rlabel viali 590 -125 615 -90 1 out
<< end >>
