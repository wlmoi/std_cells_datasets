magic
tech sky130A
timestamp 1744705058
<< locali >>
rect 2115 1045 2140 1050
rect 130 1025 465 1045
rect 130 660 155 1025
rect 1250 1020 2140 1045
rect 390 770 435 780
rect 945 775 990 785
rect 390 745 400 770
rect 425 750 465 770
rect 910 755 955 775
rect 425 745 435 750
rect 390 740 435 745
rect 945 745 955 755
rect 980 745 990 775
rect -220 640 155 660
rect -220 -440 -200 640
rect 130 590 155 640
rect 95 580 175 590
rect 95 545 115 580
rect 165 545 175 580
rect 95 535 175 545
rect 130 480 160 535
rect -125 250 -65 265
rect -125 215 -110 250
rect -75 245 -65 250
rect 270 245 330 255
rect 400 245 425 740
rect 945 735 990 745
rect 1480 675 1540 685
rect 1425 670 1540 675
rect 1425 650 1490 670
rect 1480 640 1490 650
rect 1530 640 1540 670
rect 1480 625 1540 640
rect 1500 265 1525 625
rect 2115 595 2140 1020
rect 2265 365 2335 380
rect 2265 325 2280 365
rect 2320 325 2335 365
rect 2265 310 2335 325
rect 1545 270 1600 285
rect 2280 280 2305 310
rect 1545 265 1555 270
rect 1500 245 1555 265
rect -75 225 -2 245
rect -75 215 -65 225
rect -125 200 -65 215
rect -45 -100 -25 225
rect 200 220 285 245
rect 270 215 285 220
rect 315 220 425 245
rect 1545 240 1555 245
rect 1590 265 1600 270
rect 1590 245 1625 265
rect 1590 240 1600 245
rect 475 220 975 240
rect 1545 230 1600 240
rect 2770 235 2825 245
rect 2720 230 2825 235
rect 315 215 330 220
rect 270 200 330 215
rect 145 -25 170 -7
rect 115 -35 190 -25
rect 115 -60 140 -35
rect 170 -60 190 -35
rect 115 -70 190 -60
rect 475 -100 500 220
rect 955 -65 975 220
rect 2720 215 2785 230
rect 2770 195 2785 215
rect 2815 195 2825 230
rect 2770 180 2825 195
rect 1615 150 1715 170
rect 1615 140 1635 150
rect 1315 120 1635 140
rect 1500 -65 1550 -55
rect -45 -125 500 -100
rect 945 -75 1000 -65
rect 1500 -70 1510 -65
rect 945 -100 960 -75
rect 990 -100 1000 -75
rect 1460 -90 1510 -70
rect 1500 -95 1510 -90
rect 1540 -95 1550 -65
rect 1500 -100 1550 -95
rect 945 -115 1000 -100
rect 430 -160 480 -150
rect 430 -190 440 -160
rect 470 -165 480 -160
rect 975 -165 1000 -115
rect 470 -190 500 -165
rect 945 -190 1000 -165
rect 430 -200 480 -190
rect -220 -460 495 -440
<< viali >>
rect 400 745 425 770
rect 955 745 980 775
rect 115 545 165 580
rect -110 215 -75 250
rect 1490 640 1530 670
rect 2280 325 2320 365
rect 285 215 315 245
rect 1555 240 1590 270
rect 140 -60 170 -35
rect 2785 195 2815 230
rect 960 -100 990 -75
rect 1510 -95 1540 -65
rect 440 -190 470 -160
<< metal1 >>
rect 390 770 435 780
rect 390 745 400 770
rect 425 745 435 770
rect 390 740 435 745
rect 945 775 990 785
rect 945 745 955 775
rect 980 745 990 775
rect 945 735 990 745
rect 1480 670 1540 685
rect 1480 640 1490 670
rect 1530 640 1540 670
rect 1480 625 1540 640
rect 1615 635 2305 660
rect 95 580 175 590
rect 95 545 115 580
rect 165 545 175 580
rect 95 535 175 545
rect 1615 420 1640 635
rect 1420 395 1640 420
rect 1000 310 1030 365
rect 1000 285 1060 310
rect -125 250 -65 265
rect -125 215 -110 250
rect -75 215 -65 250
rect -125 200 -65 215
rect 270 245 330 255
rect 270 215 285 245
rect 315 215 330 245
rect 1030 220 1060 285
rect 270 200 330 215
rect 420 170 745 200
rect 115 -35 190 -25
rect 420 -35 445 170
rect 1420 60 1445 395
rect 2280 380 2305 635
rect 2265 365 2335 380
rect 2265 325 2280 365
rect 2320 325 2335 365
rect 2265 310 2335 325
rect 1545 270 1600 285
rect 1545 240 1555 270
rect 1590 240 1600 270
rect 1545 230 1600 240
rect 2770 230 2825 245
rect 2770 195 2785 230
rect 2815 195 2825 230
rect 2770 180 2825 195
rect 1420 35 1540 60
rect 115 -60 140 -35
rect 170 -60 445 -35
rect 1520 -55 1540 35
rect 115 -65 445 -60
rect 1500 -65 1550 -55
rect 115 -70 190 -65
rect 945 -75 1000 -65
rect 945 -100 960 -75
rect 990 -100 1000 -75
rect 1500 -95 1510 -65
rect 1540 -95 1550 -65
rect 1500 -100 1550 -95
rect 945 -115 1000 -100
rect 430 -160 480 -150
rect 430 -190 440 -160
rect 470 -190 480 -160
rect 430 -200 480 -190
use and_common_3  and_common_3_0 /foss/designs/eda/and
timestamp 1744697173
transform 1 0 405 0 1 475
box 0 -110 1020 590
use and_common_3  and_common_3_1
timestamp 1744697173
transform 1 0 440 0 -1 110
box 0 -110 1020 590
use inv2  inv2_0 /foss/designs/eda/and
timestamp 1743223184
transform 1 0 135 0 1 328
box -140 -335 125 175
use or_common_3  or_common_3_0
timestamp 1744705058
transform 1 0 1690 0 1 110
box -65 -185 1030 485
<< labels >>
rlabel viali 285 215 315 245 1 sel_out
rlabel viali 140 -60 170 -35 1 gnd
rlabel viali 115 545 165 580 1 vdd
rlabel viali 1510 -95 1540 -65 1 out_and2
rlabel viali 440 -190 470 -160 1 in_b
rlabel viali 960 -100 990 -75 1 in2_and2
rlabel viali 955 745 980 775 1 in_a
rlabel viali -110 215 -75 250 1 in_sel
rlabel viali 1490 640 1530 670 1 out_and1
rlabel viali 1555 240 1590 270 1 in1_or
rlabel viali 2280 325 2320 365 1 in2_or
rlabel viali 2785 195 2815 230 1 out_mux
rlabel viali 400 745 425 770 1 in1_and1
<< end >>
