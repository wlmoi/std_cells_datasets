magic
tech sky130A
timestamp 1744708989
<< locali >>
rect 120 1180 530 1200
rect 120 695 145 1180
rect 1320 1170 1985 1200
rect 455 925 505 935
rect 1030 930 1090 940
rect 975 925 1090 930
rect 455 895 465 925
rect 495 905 535 925
rect 975 910 1045 925
rect 495 895 505 905
rect 455 885 505 895
rect 1030 890 1045 910
rect 1080 890 1090 925
rect -265 665 145 695
rect -265 -470 -235 665
rect 120 605 145 665
rect 105 595 185 605
rect 105 565 125 595
rect 170 565 185 595
rect 105 550 185 565
rect 135 490 155 550
rect -150 250 -85 260
rect -150 215 -135 250
rect -95 245 -85 250
rect 250 245 300 250
rect -95 215 0 245
rect 205 240 300 245
rect 470 240 490 885
rect 1030 875 1090 890
rect 1535 830 1595 840
rect 1535 825 1545 830
rect 1490 805 1545 825
rect 1535 795 1545 805
rect 1585 810 1680 830
rect 1585 795 1595 810
rect 1535 785 1595 795
rect 1465 310 1550 325
rect 1465 270 1480 310
rect 1535 270 1550 310
rect 1465 260 1550 270
rect 1655 265 1680 810
rect 1960 520 1985 1170
rect 2425 315 2505 330
rect 2425 285 2440 315
rect 2495 285 2505 315
rect 2425 275 2505 285
rect 205 225 260 240
rect 250 215 260 225
rect 290 220 490 240
rect 290 215 300 220
rect -150 205 -85 215
rect -60 -190 -30 215
rect 250 210 300 215
rect 300 160 1035 185
rect 140 -45 165 0
rect 115 -55 185 -45
rect 115 -90 125 -55
rect 175 -90 185 -55
rect 115 -100 185 -90
rect 300 -190 330 160
rect 1015 -30 1035 160
rect 1495 55 1520 260
rect 1640 240 1725 265
rect 1640 200 1665 240
rect 1705 225 1725 240
rect 1705 200 1755 225
rect 2455 210 2475 275
rect 1640 190 1755 200
rect 2430 190 2475 210
rect 2965 180 3020 195
rect 2930 160 2980 180
rect 2965 155 2980 160
rect 3005 155 3020 180
rect 2965 140 3020 155
rect 1495 25 1600 55
rect 1015 -50 1080 -30
rect -60 -215 330 -190
rect 465 -190 525 -180
rect 1060 -185 1080 -50
rect 1570 -90 1600 25
rect 1560 -100 1610 -90
rect 1560 -105 1570 -100
rect 1520 -125 1570 -105
rect 1560 -130 1570 -125
rect 1600 -130 1610 -100
rect 1560 -140 1610 -130
rect 465 -220 480 -190
rect 520 -200 525 -190
rect 1045 -195 1095 -185
rect 1045 -200 1055 -195
rect 520 -220 565 -200
rect 1005 -220 1055 -200
rect 465 -235 525 -220
rect 1045 -225 1055 -220
rect 1085 -225 1095 -195
rect 1045 -240 1095 -225
rect -265 -495 560 -470
<< viali >>
rect 465 895 495 925
rect 1045 890 1080 925
rect 125 565 170 595
rect -135 215 -95 250
rect 1545 795 1585 830
rect 1480 270 1535 310
rect 2440 285 2495 315
rect 260 215 290 240
rect 125 -90 175 -55
rect 1665 200 1705 240
rect 2980 155 3005 180
rect 1570 -130 1600 -100
rect 480 -220 520 -190
rect 1055 -225 1085 -195
<< metal1 >>
rect 455 925 505 935
rect 455 895 465 925
rect 495 895 505 925
rect 455 885 505 895
rect 1030 925 1090 940
rect 1030 890 1045 925
rect 1080 890 1090 925
rect 1030 875 1090 890
rect 1535 830 1595 840
rect 1535 795 1545 830
rect 1585 795 1595 830
rect 1535 785 1595 795
rect 105 595 185 605
rect 105 565 125 595
rect 170 565 185 595
rect 105 550 185 565
rect 1495 580 2470 600
rect -150 250 -85 260
rect -150 215 -135 250
rect -95 215 -85 250
rect -150 205 -85 215
rect 250 240 300 250
rect 250 215 260 240
rect 290 215 300 240
rect 250 210 300 215
rect 1090 185 1110 520
rect 1495 325 1525 580
rect 2445 330 2470 580
rect 1465 310 1550 325
rect 1465 270 1480 310
rect 1535 270 1550 310
rect 2425 315 2505 330
rect 2425 285 2440 315
rect 2495 285 2505 315
rect 2425 275 2505 285
rect 1465 260 1550 270
rect 1640 240 1725 265
rect 1640 200 1665 240
rect 1705 200 1725 240
rect 1640 190 1725 200
rect 2965 180 3020 195
rect 455 135 810 165
rect 1365 135 1665 165
rect 2965 155 2980 180
rect 3005 155 3020 180
rect 2965 140 3020 155
rect 115 -55 185 -45
rect 455 -55 480 135
rect 1630 130 1665 135
rect 1630 100 1850 130
rect 115 -90 125 -55
rect 175 -80 480 -55
rect 175 -90 185 -80
rect 115 -100 185 -90
rect 1560 -100 1610 -90
rect 1560 -130 1570 -100
rect 1600 -130 1610 -100
rect 1560 -140 1610 -130
rect 465 -190 525 -180
rect 465 -220 480 -190
rect 520 -220 525 -190
rect 465 -235 525 -220
rect 1045 -195 1095 -185
rect 1045 -225 1055 -195
rect 1085 -225 1095 -195
rect 1045 -240 1095 -225
use and_common_3  and_common_3_0
timestamp 1744697173
transform 1 0 473 0 1 629
box 0 -110 1020 590
use and_common_3  and_common_3_1
timestamp 1744697173
transform 1 0 502 0 -1 75
box 0 -110 1020 590
use inverter_common  inverter_common_0
timestamp 1743223184
transform 1 0 140 0 1 335
box -140 -335 125 175
use or_common_3  or_common_3_0
timestamp 1744707046
transform 1 0 1819 0 1 58
box -65 -185 1115 485
<< labels >>
rlabel viali -135 215 -95 250 1 in_sel
rlabel viali 125 565 170 595 1 vdd
rlabel viali 125 -90 175 -55 1 gnd
rlabel viali 260 215 290 240 1 out_sel
rlabel viali 465 895 495 925 1 in1_and1
rlabel viali 1045 890 1080 925 1 in_a
rlabel viali 480 -220 520 -190 1 in_b
rlabel viali 1055 -225 1085 -195 1 in2_and2
rlabel viali 1570 -130 1600 -100 1 out_and2
rlabel viali 1545 795 1585 830 1 out_and1
rlabel viali 1665 200 1705 240 1 in1_or
rlabel viali 2980 155 3005 180 1 mux_out
<< end >>
