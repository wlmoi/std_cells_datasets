magic
tech sky130A
timestamp 1744527239
<< nwell >>
rect -245 20 300 140
<< nmos >>
rect -70 -155 -50 -85
rect 180 -155 200 -85
<< pmos >>
rect -70 50 -50 115
rect 180 50 200 115
<< ndiff >>
rect -130 -100 -70 -85
rect -130 -145 -120 -100
rect -90 -145 -70 -100
rect -130 -155 -70 -145
rect -50 -100 5 -85
rect -50 -140 -30 -100
rect -5 -140 5 -100
rect -50 -155 5 -140
rect 125 -100 180 -85
rect 125 -140 135 -100
rect 160 -140 180 -100
rect 125 -155 180 -140
rect 200 -100 255 -85
rect 200 -140 220 -100
rect 245 -140 255 -100
rect 200 -155 255 -140
<< pdiff >>
rect -130 105 -70 115
rect -130 60 -120 105
rect -90 60 -70 105
rect -130 50 -70 60
rect -50 100 5 115
rect -50 65 -30 100
rect -5 65 5 100
rect -50 50 5 65
rect 125 105 180 115
rect 125 60 135 105
rect 160 60 180 105
rect 125 50 180 60
rect 200 105 255 115
rect 200 60 220 105
rect 245 60 255 105
rect 200 50 255 60
<< ndiffc >>
rect -120 -145 -90 -100
rect -30 -140 -5 -100
rect 135 -140 160 -100
rect 220 -140 245 -100
<< pdiffc >>
rect -120 60 -90 105
rect -30 65 -5 100
rect 135 60 160 105
rect 220 60 245 105
<< psubdiff >>
rect -220 -105 -165 -85
rect -220 -140 -205 -105
rect -180 -140 -165 -105
rect -220 -155 -165 -140
rect 295 -100 345 -85
rect 295 -140 305 -100
rect 335 -140 345 -100
rect 295 -155 345 -140
<< nsubdiff >>
rect -220 100 -165 115
rect -220 65 -205 100
rect -180 65 -165 100
rect -220 50 -165 65
<< psubdiffcont >>
rect -205 -140 -180 -105
rect 305 -140 335 -100
<< nsubdiffcont >>
rect -205 65 -180 100
<< poly >>
rect -70 115 -50 130
rect 180 115 200 130
rect -70 -5 -50 50
rect -110 -15 -50 -5
rect -110 -40 -105 -15
rect -75 -40 -50 -15
rect -110 -50 -50 -40
rect -70 -85 -50 -50
rect 180 -5 200 50
rect 180 -15 245 -5
rect 180 -40 210 -15
rect 235 -40 245 -15
rect 180 -50 245 -40
rect 180 -85 200 -50
rect -70 -170 -50 -155
rect 180 -170 200 -155
<< polycont >>
rect -105 -40 -75 -15
rect 210 -40 235 -15
<< locali >>
rect -30 175 245 195
rect -30 115 -5 175
rect 225 115 245 175
rect -220 100 -165 115
rect -220 65 -205 100
rect -180 95 -165 100
rect -130 105 -80 115
rect -130 95 -120 105
rect -180 75 -120 95
rect -180 65 -165 75
rect -220 50 -165 65
rect -130 60 -120 75
rect -90 60 -80 105
rect -130 50 -80 60
rect -40 100 5 115
rect -40 65 -30 100
rect -5 65 5 100
rect -40 50 5 65
rect 125 105 170 115
rect 125 60 135 105
rect 160 60 170 105
rect 125 50 170 60
rect 210 105 255 115
rect 210 60 220 105
rect 245 60 255 105
rect 210 50 255 60
rect 135 -5 160 50
rect -110 -15 -70 -5
rect -110 -40 -105 -15
rect -75 -40 -70 -15
rect -110 -50 -70 -40
rect -30 -10 160 -5
rect -30 -45 35 -10
rect 85 -45 160 -10
rect -30 -50 160 -45
rect 200 -15 245 -5
rect 200 -40 210 -15
rect 235 -40 245 -15
rect 200 -50 245 -40
rect -30 -85 -5 -50
rect -220 -105 -165 -85
rect -220 -140 -205 -105
rect -180 -110 -165 -105
rect -130 -100 -80 -85
rect -130 -110 -120 -100
rect -180 -135 -120 -110
rect -180 -140 -165 -135
rect -220 -155 -165 -140
rect -130 -145 -120 -135
rect -90 -145 -80 -100
rect -130 -155 -80 -145
rect -40 -100 5 -85
rect -40 -140 -30 -100
rect -5 -140 5 -100
rect -40 -155 5 -140
rect 45 -225 65 -50
rect 135 -85 160 -50
rect 125 -100 170 -85
rect 125 -140 135 -100
rect 160 -140 170 -100
rect 125 -155 170 -140
rect 210 -100 255 -85
rect 210 -140 220 -100
rect 245 -110 255 -100
rect 295 -100 345 -85
rect 295 -110 305 -100
rect 245 -130 305 -110
rect 245 -140 255 -130
rect 210 -155 255 -140
rect 295 -140 305 -130
rect 335 -140 345 -100
rect 295 -155 345 -140
rect 455 -225 475 -50
rect 45 -245 475 -225
<< viali >>
rect -205 65 -180 100
rect 35 -45 85 -10
rect -205 -140 -180 -105
rect 305 -140 335 -100
<< metal1 >>
rect -220 100 -165 115
rect -220 65 -205 100
rect -180 65 -165 100
rect -220 50 -165 65
rect -30 -10 160 -5
rect -30 -45 35 -10
rect 85 -45 160 -10
rect -30 -50 160 -45
rect -220 -105 -165 -85
rect -220 -140 -205 -105
rect -180 -140 -165 -105
rect -220 -155 -165 -140
rect 295 -100 345 -85
rect 295 -140 305 -100
rect 335 -140 345 -100
rect 295 -155 345 -140
use inv2  inv2_0 /foss/designs/eda/inverter
timestamp 1743223184
transform 1 0 580 0 1 80
box -140 -335 125 175
<< labels >>
rlabel nwell -205 65 -180 100 1 vdd
rlabel polycont -105 -40 -75 -15 1 in1
rlabel viali 35 -45 85 -10 1 out
rlabel polycont 210 -40 235 -15 1 in2
rlabel metal1 -205 -140 -180 -105 1 gnd
rlabel metal1 305 -140 335 -100 1 gnd
rlabel space 580 -240 605 -220 1 gnd
rlabel space 565 190 605 220 1 vdd
rlabel space 610 -35 635 -10 1 out
<< end >>
