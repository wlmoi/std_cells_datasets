magic
tech sky130A
timestamp 1744697173
<< locali >>
rect 415 575 490 590
rect 415 570 435 575
rect 55 550 435 570
rect 55 415 75 550
rect 415 545 435 550
rect 475 570 490 575
rect 475 550 850 570
rect 475 545 490 550
rect 415 535 490 545
rect 825 450 850 550
rect 60 300 110 305
rect 455 300 505 310
rect 60 275 70 300
rect 100 295 110 300
rect 100 275 140 295
rect 415 280 465 300
rect 60 265 110 275
rect 455 270 465 280
rect 495 270 505 300
rect 455 260 505 270
rect 965 200 1020 210
rect 900 180 975 200
rect 965 175 975 180
rect 1010 175 1020 200
rect 965 165 1020 175
rect 570 -65 640 -50
rect 570 -95 590 -65
rect 625 -95 640 -65
rect 570 -110 640 -95
<< viali >>
rect 435 545 475 575
rect 70 275 100 300
rect 465 270 495 300
rect 710 180 735 205
rect 975 175 1010 200
rect 590 -95 625 -65
<< metal1 >>
rect 415 575 490 590
rect 415 545 435 575
rect 475 545 490 575
rect 415 535 490 545
rect 265 480 725 500
rect 265 310 285 480
rect 60 300 110 305
rect 60 275 70 300
rect 100 275 110 300
rect 60 265 110 275
rect 455 300 505 310
rect 455 270 465 300
rect 495 270 505 300
rect 455 260 505 270
rect 700 220 725 480
rect 695 205 750 220
rect 695 180 710 205
rect 735 180 750 205
rect 695 165 750 180
rect 965 200 1020 210
rect 965 175 975 200
rect 1010 175 1020 200
rect 965 165 1020 175
rect 305 -65 330 70
rect 570 -65 640 -50
rect 835 -65 865 -40
rect 305 -90 590 -65
rect 570 -95 590 -90
rect 625 -90 865 -65
rect 625 -95 640 -90
rect 570 -110 640 -95
use inv2  inv2_0
timestamp 1743223184
transform 1 0 835 0 1 295
box -140 -335 125 175
use nand  nand_0 /foss/designs/eda/nand
timestamp 1744185391
transform 1 0 225 0 1 345
box -225 -345 315 105
<< labels >>
rlabel viali 435 545 475 575 1 vdd
rlabel viali 465 270 495 300 1 in2
rlabel viali 70 275 100 300 1 in1
rlabel viali 590 -95 625 -65 1 gnd
rlabel viali 975 175 1010 200 1 out
<< end >>
