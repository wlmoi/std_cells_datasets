magic
tech sky130A
timestamp 1744815696
<< locali >>
rect 2090 965 2545 1000
rect 4620 985 4695 1000
rect 4620 980 4635 985
rect 4485 960 4635 980
rect 4620 955 4635 960
rect 4680 955 4695 985
rect 4620 940 4695 955
rect -155 795 -65 815
rect -155 745 -135 795
rect -85 790 -65 795
rect -85 755 5 790
rect -85 745 -65 755
rect -155 725 -65 745
rect -345 545 310 580
rect -345 -490 -315 545
rect 4320 505 4345 535
rect 4320 495 4390 505
rect 4320 470 4335 495
rect 4375 470 4390 495
rect 4320 455 4390 470
rect 2355 255 2470 270
rect 2355 210 2375 255
rect 2450 210 2470 255
rect 2355 190 2470 210
rect -195 -205 -120 -190
rect -195 -240 -180 -205
rect -135 -215 -120 -205
rect 395 -200 425 55
rect 2235 -200 2240 -195
rect 395 -215 2240 -200
rect 2790 -210 2810 35
rect -135 -240 -55 -215
rect 150 -230 2240 -215
rect 2440 -230 2810 -210
rect 150 -235 2235 -230
rect -195 -260 -120 -240
rect 75 -485 110 -450
rect 930 -465 1075 -440
rect 930 -485 960 -465
rect 75 -490 960 -485
rect -345 -525 960 -490
rect 1050 -485 1075 -465
rect 2375 -485 2410 -455
rect 1050 -525 2410 -485
rect 930 -555 1075 -525
<< viali >>
rect 4635 955 4680 985
rect -135 745 -85 795
rect 4335 470 4375 495
rect 2375 210 2450 255
rect -180 -240 -135 -205
rect 960 -525 1050 -465
<< metal1 >>
rect 4620 985 4695 1000
rect 4620 955 4635 985
rect 4680 955 4695 985
rect 4620 940 4695 955
rect -155 795 -65 815
rect -155 745 -135 795
rect -85 745 -65 795
rect -155 725 -65 745
rect 4320 495 4390 505
rect 4320 470 4335 495
rect 4375 470 4390 495
rect 4320 455 4390 470
rect 2355 255 2470 270
rect 90 220 715 255
rect 2180 220 2375 255
rect 90 30 130 220
rect 2355 210 2375 220
rect 2450 215 3105 255
rect 2450 210 2470 215
rect 2355 190 2470 210
rect 2390 30 2430 190
rect -195 -205 -120 -190
rect -195 -240 -180 -205
rect -135 -240 -120 -205
rect -195 -260 -120 -240
rect 930 -465 1075 -435
rect 930 -525 960 -465
rect 1050 -525 1075 -465
rect 930 -555 1075 -525
use ff_common  ff_common_0
timestamp 1744728648
transform 1 0 210 0 1 535
box -210 -535 1975 825
use ff_common  ff_common_1
timestamp 1744728648
transform 1 0 2604 0 1 517
box -210 -535 1975 825
use inverter_common  inverter_common_0
timestamp 1743223184
transform 1 0 2375 0 1 -120
box -140 -335 125 175
use inverter_common  inverter_common_1
timestamp 1743223184
transform 1 0 85 0 1 -125
box -140 -335 125 175
<< labels >>
rlabel viali -180 -240 -135 -205 1 in_clk
rlabel viali 2375 210 2450 255 1 vdd
rlabel viali -135 745 -85 795 1 in_d
rlabel viali 960 -525 1050 -465 1 gnd
rlabel viali 4635 955 4680 985 1 out_q
rlabel viali 4335 470 4375 495 1 out_q_not
<< end >>
